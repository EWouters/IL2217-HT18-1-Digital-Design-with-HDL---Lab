--USE WORK.ALL;
--USE WORK.package_MicroAssemblyCode.ALL;
--
--LIBRARY IEEE;
--USE IEEE.std_logic_1164.all;
--USE IEEE.std_logic_signed.all;
--
--ENTITY videoComposer_fpga IS
--	GENERIC (
--		Size  : INTEGER:=8; -- # bits in word
--		ASize : INTEGER:=3  -- # bits in address
--	);
--	PORT (
--		Clk   : IN STD_LOGIC;
--		Reset : IN STD_LOGIC;
--		Ready : OUT STD_LOGIC;
--		q     : OUT STD_LOGIC_VECTOR(7 downto 0)
--	);
--END videoComposer_fpga;
--
--ARCHITECTURE behaviour OF videoComposer_fpga IS
----	CONSTANT ROM : Program_Type := (
--	--| IE | Dest | Src1 | Src2 | OpAlu | OpShift | OE |
----	( ...
----	);
--	COMPONENT dataPath
--		GENERIC (
--			Size  : INTEGER := 8; -- # bits in word
--			ASize : INTEGER := 3  -- # bits in address
--		);
--		PORT (
--			InPort  : IN STD_LOGIC_VECTOR(Size-1 DOWNTO 0);
--			OutPort : OUT STD_LOGIC_VECTOR(Size-1 DOWNTO 0);
--			Clk     : IN STD_LOGIC;
--			Instr   : IN Instruction_Type
--		);
--	END COMPONENT;
--	
--	COMPONENT single_port_ram
----		PORT
----		(
----		...
----		);
--	END COMPONENT;
--	
--	COMPONENT single_port_rom
----		PORT
----		(
----		...
----		);
--	END COMPONENT;
--	
--	-- Datapath signals
--	SIGNAL in_port : STD_LOGIC_VECTOR(Size-1 DOWNTO 0);
--	SIGNAL out_port : STD_LOGIC_VECTOR(Size-1 DOWNTO 0);
--	SIGNAL instr : Instruction_type := ( '0' , Rx , Rx , Rx , OpX , OpX , '0' );
--	
--	TYPE State_Type IS (reset_state,S_ReadRed, S_ReadGreenWriteRed, S_ReadBlueWriteGreen,
--		S_ProcessBlue, S_WriteBlue, S_Idle);
--	
--	SIGNAL current_state, next_state : State_Type;
--		-- Instr counter for the datapath
--	SIGNAL current_counter, next_counter : INTEGER := 0;
--	
--	SIGNAL read_address,next_read_address,write_address,next_write_address:
--		STD_LOGIC_VECTOR(?? DOWNTO 0);
--	
--	SIGNAL read_data,write_data_out:STD_LOGIC_VECTOR(7 downto 0);
--	SIGNAL wr_en,wr_ram:STD_LOGIC:='0';
--	
--BEGIN
--	instr <= ROM(current_counter);
--	in_port <= read_data;
--	
--	COMB: PROCESS(current_state, current_counter, read_address, write_address,
--		read_data,out_port)
--	BEGIN
--		next_state <= current_state;
--		next_counter <= current_counter;
--		Ready <= '0';
--		next_read_address<=(others=>'0');
--		next_write_address<=(others=>'0');
--		wr_en<='0';
--		CASE current_state IS
--			WHEN reset_state =>
--				next_read_address<=(others=>'0');
--				next_write_address<=(others=>'0');
--				wr_en<='0';
--				next_state<=S_ReadRed;
--				next_counter <= 0;
--			WHEN S_ReadRed => -- ROM Instr 0
--				next_state<=S_ReadGreenWriteRed;
--				next_counter <= 1;
--				next_read_address<=read_address+1;
--			WHEN S_ReadGreenWriteRed => -- ROM Instr 1
--				wr_en<='1';
--				next_counter <= 2;
--				next_state <= S_ReadBlueWriteGreen;
--				next_read_address<=read_address+1;
--				next_write_address<=write_address+1;
--			WHEN S_ReadBlueWriteGreen => -- ROM Instr 2
--				wr_en<='1';
--				next_counter <= 3;
--				next_state <= S_ProcessBlue;
--				next_read_address<=read_address+1;
--				next_write_address<=write_address+1;
--			WHEN S_ProcessBlue => -- ROM Instr 3-8
--				IF current_counter < 9 THEN
--					next_counter <= current_counter + 1;
--					next_state <= S_ProcessBlue;
--				ELSE
--					IF out_port = "00000000" THEN
--						next_counter <= 10;
--					ELSE
--						next_counter <= 11;
--					END IF;
--					next_state <= S_WriteBlue;
--				END IF;
--			WHEN S_WriteBlue => -- ROM Instr 10 or 11
--				wr_en<='1';
--				next_write_address<=write_address+1;
--				next_state <= S_Idle;
--			WHEN S_Idle =>
--				if (read_address=57600) then
--					Ready <= '1';
--				else
--					next_state<=S_ReadRed;
--					next_counter<=0;
--				end if;
--			WHEN OTHERS =>
--				ASSERT false
--				report "illegal FSM state, testbench error"
--				severity error;
--		END CASE;
--	END PROCESS;
--	
--	P_SYNCH: PROCESS(Clk,reset)
--	BEGIN
--		IF (reset='0') then
--			current_state<=reset_state;
--			current_counter<=0;
--		ELSIF Clk'EVENT AND Clk = '1' THEN
--			read_address <= next_read_address;
--			write_address <= next_write_address;
--			current_state <= next_state;
--			current_counter <= next_counter;
--		END IF;
--	END PROCESS;
--	
--	U_dataPath : dataPath
--		GENERIC MAP(Size => Size, ASize => ASize)
--		PORT MAP( InPort => in_port,
--			OutPort => out_port,
--			Clk => Clk,
--			Instr => instr
--		);
--	
--	Read_ROM:single_port_rom port map (read_address,read_data);
--	
--	Write_RAM:single_port_ram port map (write_address,wr_ram,out_port,q);
--	
--	-- Ensure a late cycle write to allow address to change first 
--	wr_ram<=wr_en AND not(clk);
--
--END behaviour;